library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity P3 is
port(

input : std_logic

);
end P3;



architecture first of P3 is

begin

test1 : block
begin

end block test1;





end first;