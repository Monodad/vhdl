library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.itc.all;
use work.itc_lcd.all;

entity gen_font is
	port (
		x                                                    : in integer range 0 to 127;
		y                                                       : in integer range 0 to 159;
		font_start                                              : in std_logic;
		font_busy                                               : out std_logic;
		clk, rst_n                                              : in std_logic;
		data                                                    : in string(1 to 5);
		text_color                                              : in l_px_t;
		bg_color                                                : in l_px_t;
		clear                                                   : in std_logic;
		lcd_sclk, lcd_mosi, lcd_ss_n, lcd_dc, lcd_bl, lcd_rst_n : out std_logic
	);
end gen_font;

architecture arch of gen_font is
	signal start_draw : std_logic;
	signal l_addr, l_addr_p, addr : l_addr_t;
	signal l_data : l_px_t;
	signal wr_ena : std_logic;
	signal q : std_logic_vector(0 downto 0);
	type status_t is (idle, draw, clear_screen);
	signal status : status_t;
	signal p_count : integer range 0 to 20;
	signal data_y, data_x : integer range 0 to 20;
	signal lcd_x : integer range 0 to 127;
	signal lcd_y : integer range 0 to 159;
	signal first_px : l_addr_t;
	signal count : integer range 0 to 10;
	signal l_clear : std_logic;
begin
	edge_inst : entity work.edge(arch)
		port map(
			clk     => clk,
			rst_n   => rst_n,
			sig_in  => font_start,
			rising  => start_draw,
			falling => open
		);
	edge_inst1 : entity work.edge(arch)
		port map(
			clk     => clk,
			rst_n   => rst_n,
			sig_in  => clear,
			rising  => l_clear,
			falling => open
		);
	lcd_inst : entity work.lcd(arch)
		port map(
			clk        => clk,
			rst_n      => rst_n,
			lcd_sclk   => lcd_sclk,
			lcd_mosi   => lcd_mosi,
			lcd_ss_n   => lcd_ss_n,
			lcd_dc     => lcd_dc,
			lcd_bl     => lcd_bl,
			lcd_rst_n  => lcd_rst_n,
			brightness => 100,
			wr_ena     => wr_ena,
			addr       => l_addr,
			data       => l_data
		);
	font_inst : entity work.Font(SYN)
		port map(
			address => std_logic_vector(to_unsigned(l_addr_p, 15)),
			clock   => clk,
			q       => q
		);
	l_data <= x"000000" when (q = "1") and (status /= clear_screen) else
		bg_color when status = clear_screen else x"26B2E3";
	process (clk, rst_n)
	begin
		if (rst_n = '0') then
			wr_ena <= '0';
			status <= clear_screen;
			count <= 0;
			data_x <= 0;
			data_y <= 0;
			count <= 0;
			addr <= 0;
		elsif rising_edge(clk) then
			case status is
				when idle =>
					if (start_draw = '1') then
						p_count <= data'length;
						status <= draw;
						wr_ena <= '1';
						font_busy <= '1';
						--lcd_x <= x;
						lcd_y <= y;
					else
						wr_ena <= '0';
						font_busy <= '0';
					end if;
					if (l_clear = '1') then
						wr_ena <= '1';
						font_busy <= '1';
						addr <= 0;
						status <= clear_screen;
					else
						wr_ena <= '0';
						font_busy <= '0';
					end if;
				when draw =>
					if (data_x = 10) then
						data_y <= data_y + 1;
						data_x <= 0;
					else
						data_x <= data_x + 1;
					end if;
					if (data_y = 20) then
						data_y <= 0;

						if (count = data'length) then
							status <= idle;
							count <= 0;
							data_x <= 0;
							data_y <= 0;
							font_busy <= '1';
						else
							count <= count + 1;
						end if;
					end if;
					if (((data_x) > 127) or ((data_y + y) > 159)) then
						wr_ena <= '0';
					else
						wr_ena <= '1';
					end if;
				when clear_screen =>
					if (addr = addr'high) then
						addr <= 0;
						status <= idle;
					else
						addr <= addr + 1;
					end if;
				when others =>
					status <= idle;
			end case;

		end if;
	end process;
	l_addr_p <= 950 * data_y + data_x + first_px;
	first_px <= (character'pos(data(count + 1)) - 32) * 10;
	l_addr <= 128 * (data_y + y) + data_x + (count * 11) when status /= clear_screen else addr;
end arch;
